module image_bank
#(  
    parameter HEX_IDX = 3,
    parameter LOAD_MEM = 0
)
(
    input logic clk,
    input logic rst_n,
    input logic [6:0] raddr,
    input logic [6:0] waddr,
    input logic re,
    input logic we,
    input logic [3071:0] wdata,
    input logic [1:0] idx,
    output logic [3071:0] rdata
);

    // Image bank
    (* ramstyle = "mlab" *) logic [3071:0] bank [0:63];
    // logic [3071:0] bank [0:85];

    // Write enable
    always_ff @(posedge clk) begin
        if (we) begin
            bank[waddr] <= wdata;
        end
    end

    // Read enable
    always_ff @(posedge clk, negedge rst_n) begin
        if (~rst_n) begin
            rdata <= '0;
        end
        else
        if (re) begin
            rdata <= bank[raddr];
        end
    end

    // Load test.hex to image bank for testing purpose
    initial begin
        if (LOAD_MEM == 1)
            if (HEX_IDX == 0)
                $readmemh("I:/ECE554/Testing/Bank0.hex", bank);
            else if (HEX_IDX == 1)
                $readmemh("I:/ECE554/Testing/Bank1.hex", bank);
            else if (HEX_IDX == 2)
                $readmemh("I:/ECE554/Testing/Bank2.hex", bank);
        // if (LOAD_MEM == 1)
        //     if (HEX_IDX == 0)
        //         $readmemh("C:\\Users\\asus\\Desktop\\ECE554\\ECE554\-SP24\\Final_Project\\RTL\\coproc\\Bank0.hex", bank);
        //     else if (HEX_IDX == 1)
        //         $readmemh("C:\\Users\\asus\\Desktop\\ECE554\\ECE554\-SP24\\Final_Project\\RTL\\coproc\\Bank1.hex", bank);
        //     else if (HEX_IDX == 2)
        //         $readmemh("C:\\Users\\asus\\Desktop\\ECE554\\ECE554\-SP24\\Final_Project\\RTL\\coproc\\Bank2.hex", bank);
    end

endmodule