module pixel_sel_tb();

    // DUT Signals
    logic [3071:0] rdata0_in, rdata1_in, rdata2_in;
    logic [7:0] col_cnt;
    logic [2:0] row_sel_onehot;
    logic [35:0] rdata0_out, rdata1_out, rdata2_out;

    // Instantiate pixel select module
    pixel_sel iPexel_Sel(
        .rdata0_in(rdata0_in), .rdata1_in(rdata1_in), .rdata2_in(rdata2_in),
        .col_cnt(col_cnt), .row_sel_onehot(row_sel_onehot),
        .rdata0_out(rdata0_out), .rdata1_out(rdata1_out), .rdata2_out(rdata2_out));

    logic clk, rst_n;

    always_ff @(negedge clk, negedge rst_n) begin
        if(~rst_n)
            col_cnt <= '0;
        else
            col_cnt <= col_cnt + 1;
    end

    always_ff @(posedge clk, negedge rst_n) begin
        // TODO: to be tested, need to think about initial value
        if (~rst_n) begin
            row_sel_onehot <= 3'b001;
        end
        else if (~(|col_cnt)) begin
            row_sel_onehot <= {row_sel_onehot[1:0], row_sel_onehot[2]};
        end
    end

    initial begin
        clk = 0;
        rst_n = 0;
        rdata0_in = 3072'h00000100200300400500600700800900a00b00c00d00e00f01001101201301401501601701801901a01b01c01d01e01f02002102202302402502602702802902a02b02c02d02e02f03003103203303403503603703803903a03b03c03d03e03f04004104204304404504604704804904a04b04c04d04e04f05005105205305405505605705805905a05b05c05d05e05f06006106206306406506606706806906a06b06c06d06e06f07007107207307407507607707807907a07b07c07d07e07f08008108208308408508608708808908a08b08c08d08e08f09009109209309409509609709809909a09b09c09d09e09f0a00a10a20a30a40a50a60a70a80a90aa0ab0ac0ad0ae0af0b00b10b20b30b40b50b60b70b80b90ba0bb0bc0bd0be0bf0c00c10c20c30c40c50c60c70c80c90ca0cb0cc0cd0ce0cf0d00d10d20d30d40d50d60d70d80d90da0db0dc0dd0de0df0e00e10e20e30e40e50e60e70e80e90ea0eb0ec0ed0ee0ef0f00f10f20f30f40f50f60f70f80f90fa0fb0fc0fd0fe0ff;
        rdata1_in = 3072'h10010110210310410510610710810910a10b10c10d10e10f11011111211311411511611711811911a11b11c11d11e11f12012112212312412512612712812912a12b12c12d12e12f13013113213313413513613713813913a13b13c13d13e13f14014114214314414514614714814914a14b14c14d14e14f15015115215315415515615715815915a15b15c15d15e15f16016116216316416516616716816916a16b16c16d16e16f17017117217317417517617717817917a17b17c17d17e17f18018118218318418518618718818918a18b18c18d18e18f19019119219319419519619719819919a19b19c19d19e19f1a01a11a21a31a41a51a61a71a81a91aa1ab1ac1ad1ae1af1b01b11b21b31b41b51b61b71b81b91ba1bb1bc1bd1be1bf1c01c11c21c31c41c51c61c71c81c91ca1cb1cc1cd1ce1cf1d01d11d21d31d41d51d61d71d81d91da1db1dc1dd1de1df1e01e11e21e31e41e51e61e71e81e91ea1eb1ec1ed1ee1ef1f01f11f21f31f41f51f61f71f81f91fa1fb1fc1fd1fe1ff;
        rdata2_in = 3072'h20020120220320420520620720820920a20b20c20d20e20f21021121221321421521621721821921a21b21c21d21e21f22022122222322422522622722822922a22b22c22d22e22f23023123223323423523623723823923a23b23c23d23e23f24024124224324424524624724824924a24b24c24d24e24f25025125225325425525625725825925a25b25c25d25e25f26026126226326426526626726826926a26b26c26d26e26f27027127227327427527627727827927a27b27c27d27e27f28028128228328428528628728828928a28b28c28d28e28f29029129229329429529629729829929a29b29c29d29e29f2a02a12a22a32a42a52a62a72a82a92aa2ab2ac2ad2ae2af2b02b12b22b32b42b52b62b72b82b92ba2bb2bc2bd2be2bf2c02c12c22c32c42c52c62c72c82c92ca2cb2cc2cd2ce2cf2d02d12d22d32d42d52d62d72d82d92da2db2dc2dd2de2df2e02e12e22e32e42e52e62e72e82e92ea2eb2ec2ed2ee2ef2f02f12f22f32f42f52f62f72f82f92fa2fb2fc2fd2fe2ff;


        @(negedge clk);
        rst_n = 1;

        repeat(300) @(negedge clk);

        $stop();
    end

    always #5 clk = ~clk;

endmodule